/*
* @File name: issue_buffer
* @Author: Ruige Lee
* @Email: wut.ruigeli@gmail.com
* @Date:   2020-10-27 18:04:15
* @Last Modified by:   Ruige Lee
* @Last Modified time: 2020-10-27 18:05:43
*/

module issue_buffer #
(
	parameter DW = 100,
	parameter DP = 8,
)


(




	input CLK,
	input RSTn
	
);

endmodule








