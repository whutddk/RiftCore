
`timescale 1 ns / 1 ps





