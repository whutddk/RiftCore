/*
* @File name: writeBack
* @Author: Ruige Lee
* @Email: wut.ruigeli@gmail.com
* @Date:   2020-09-11 15:41:38
* @Last Modified by:   Ruige Lee
* @Last Modified time: 2020-10-26 17:44:45
*/

module writeBack (

	output [32*RNDEPTH-1 : 0] writeBackBuffer_qout,

	input [32*RNDEPTH-1 : 0] instr_issue,

	input [32*RNDEPTH-1 : 0] instr_commit


	
);













endmodule

