/*
* @File name: instr_fetch
* @Author: Ruige Lee
* @Email: wut.ruigeli@gmail.com
* @Date:   2020-09-11 15:40:23
* @Last Modified by:   Ruige Lee
* @Last Modified time: 2020-10-30 17:24:58
*/

module instr_fetch (
	
);


$warning("预留一拍做后处理");







endmodule


