/*
* @File name: execute
* @Author: Ruige Lee
* @Email: wut.ruigeli@gmail.com
* @Date:   2020-09-11 15:40:54
* @Last Modified by:   Ruige Lee
* @Last Modified time: 2020-09-19 15:30:42
*/

module execute (
	



);



alu i_alu();

blu i_blu();














endmodule


