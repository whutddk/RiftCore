/*
* @File name: inOrder_fifo
* @Author: Ruige Lee
* @Email: wut.ruigeli@gmail.com
* @Date:   2020-10-23 17:41:48
* @Last Modified by:   Ruige Lee
* @Last Modified time: 2020-10-23 17:58:17
*/


module inOrder_fifo (



	
	input CLK,
	input RSTn
	
);

endmodule











