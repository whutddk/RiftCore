/*
* @File name: commit
* @Author: Ruige Lee
* @Email: wut.ruigeli@gmail.com
* @Date:   2020-09-11 15:41:55
* @Last Modified by:   Ruige Lee
* @Last Modified time: 2020-10-20 17:45:29
*/

module commit (

);








//代表架构寄存器，指向128个寄存器中的地址，完成commit
wire [6*31:0] arch_x;










endmodule


