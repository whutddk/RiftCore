/*
* @File name: pc_generate
* @Author: Ruige Lee
* @Email: wut.ruigeli@gmail.com
* @Date:   2020-10-13 16:56:39
* @Last Modified by:   Ruige Lee
* @Last Modified time: 2020-10-18 15:50:41
*/

//产生的pc不是执行pc，每条指令应该对应一个pc



module pc_generate (

	input [63:0] decode_pc,



	input [63:0] blu_pc,
	input [63:0] blu_res,



	output [63:0] fetch_pc
);











































endmodule










