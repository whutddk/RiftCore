/*
* @File name: fetch
* @Author: Ruige Lee
* @Email: wut.ruigeli@gmail.com
* @Date:   2020-09-11 15:40:23
* @Last Modified by:   Ruige Lee
* @Last Modified time: 2020-09-11 15:41:13
*/

module fetch (
	
);

endmodule


