/*
* @File name: oth_issue
* @Author: Ruige Lee
* @Email: wut.ruigeli@gmail.com
* @Date:   2020-10-27 10:52:23
* @Last Modified by:   Ruige Lee
* @Last Modified time: 2020-10-27 10:52:39
*/

module oth_issue (





	input oth_issue_vaild,
	output oth_issue_ready,
	input [:] oth_issue_info,














);



















endmodule












